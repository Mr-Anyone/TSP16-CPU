`define A_TYPE 2'b00
`define M_TYPE 2'b01
`define R_TYPE 2'b10
`define B_TYPE 2'b11

`define ADD 5'b00000
`define EQUAL 5'b00001
`define OR 5'b00010
`define AND 5'b00011
`define MINUS 5'b00100

